module font_rom   (input        [4:0]   wordkey,
						 output logic [143:0] outputWord);
	always_comb
	begin
		unique case (wordkey)
			5'b00000: outputWord = 144'b000000000000011111111110011111111110011000000110011000000110011000000110011000000110011000000110011000000110011111111110011111111110000000000000; //o
												 
			5'b00001: outputWord = 144'b000000000000011000000110011000000110011000000110011000000110011111111110011111111110011000000110011000000110011000000110011000000110000000000000; //H
			
												 
			5'b00010: outputWord = 144'b000000000000001111111100001111111100000001100000000001100000000001100000000001100000000001100000000001100000001111111100001111111100000000000000; //I
												 
			5'b00011: outputWord = 144'b000000000000000111111000001111111100001100000000001100000000001100011110001100011110001100000110001100000110001111111110000111111100000000000000; //G
												 
			5'b00100: outputWord = 144'b000000000000001100000000001100000000001100000000001100000000001100000000001100000000001100000000001100000000001111111110000111111100000000000000; //L
												 
			5'b00101: outputWord = 144'b000000000000011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011011110110001110011100000000000000; //W
												 
			5'b00110: outputWord = 144'b000000000000001111111100001111111100001100000000001100000000001111111100001111111100001100000000001100000000001111111100001111111100000000000000; //E
												 
			5'b00111: outputWord = 144'b000000000000001111111110001111111110001100000000001100000000001100000000001100000000001100000000001100000000001111111110001111111110000000000000; //C
												 
			5'b01000: outputWord = 144'b000000000000000111111100001111111110001100000110001100000110001111111110001111111100001100000000001100000000001100000000001100000000000000000000; //P
			
			5'b01001: outputWord = 144'b000000000000011111111110011111111110000001100000000001100000000001100000000001100000000001100000000001100000000001100000000001100000000000000000; //T
												 
			5'b01010: outputWord = 144'b000000000000011111111110011111111110011000000000011000000000011111111110011111111110011000000000011000000000011000000000011000000000000000000000; //F
			
			5'b01011: outputWord = 144'b000001100000000011110000000111111000001111111100011111111110000001100000000001100000000001100000000001100000000001100000000001100000000000000000; //uparrow
			
			5'b01100: outputWord = 144'b000000000000000001100000000001100000000001100000000001100000000001100000000001100000011111111110001111111100000111111000000011110000000001100000; //downarrow

			default : outputWord = 144'b0; 
		endcase
	end
	
endmodule
